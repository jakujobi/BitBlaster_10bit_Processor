// Authors: John Akujobi
// Date: November, Fall, 2023
// Name: Input Logic
// Filename: inputlogic.sv
// Description: The input logic module manages external inputs to the processor.
// It includes debouncing logic for stable input signals and routes external
// data to the processor's internal bus. It plays a vital role in interfacing
// the processor with external sources like switches and buttons.

module inputlogic (
    input logic [9:0] RawData,
    input logic Peek_key,
    input logic CLK_50MHz,
    input logic RawCLK,
    input Extrn_Enable,

    output logic [9:0] databus,
    output logic [1:0] data2bit,
    output logic CLKb,
    output logic PeeKb
);

//assign databus = 10'bz;

//Debounce the keys__________________________________________
debouncer peek_debouncer (
    .A_noisy(Peek_key),
    .CLK50M(CLK_50MHz),
    .A(PeeKb)
);

debouncer clk_debouncer (
    .A_noisy(RawCLK),
    .CLK50M(CLK_50MHz),
    .A(CLKb)
);

//splice the lowest 2 bits
assign data2bit = RawData[1:0];

// //if extrn is enabled, assign raw data to databus
// assign databus = Extrn_Enable ? RawData : z;

//always comp block that assigns the data to the databus
always_comb begin
    if (Extrn_Enable) begin
        databus = RawData;
    end
    else begin
        databus = 10'bz;
    end
end

// extrn external_data_receiver (
//     .raw_data(raw_data),
//     .extrn_enable (extrn_enable),
//     .PKb(PKb)
// );


endmodule