module controller(
    input logic [9:0] INST,
    input logic [1:0] T,

    output logic [9:0] IMM,
    output logic [1:0] Rin,
    output logic [1:0] Rout,
    output logic ENW,
    output logic ENR,
    output logic Ain,
    output logic Gin,
    output logic Gout,
    output logic [3:0] ALUcont,
    output logic Ext,
    output logic IRin,
    output logic Clr
);



endmodule