module extrn (
    input logic [9:0] raw_data,
    input logic extrn_enable,

    output logic [1:0] data2,
    output logic [9:0] outdata
);


endmodule