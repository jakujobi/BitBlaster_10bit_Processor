module outputlogic(
    input logic [9:0] BUS,
    input logic [9:0] REG,
    input logic [1:0] TIME,
    input logic DONE,
    input logic Pkb,

    output logic [9:0] LED_B,
    output logic [6:0] DHEX0,
    output logic [6:0] DHEX1
    output logic [6:0] DHEX2,
    output logic [6:0] THEX,
    output logic LED_D
);





endmodule