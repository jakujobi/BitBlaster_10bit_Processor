module registerFile (
    input logic [9:0] D ,
    input logic ENW , ENR0 , ENR1 , CLKb ,
    input logic [1:0] WRA , RDA0 , RDA1 ,
    output logic [9:0] Q0 , Q1
);




endmodule