module inputlogic (

);


endmodule